interface intf(input logic clk);

endinterface